-- DTH11 controller wrapper, standalone version

library ieee;
use ieee.std_logic_1164.all;

entity dht11_sa is
	generic(
		freq:    positive range 1 to 1000 -- Clock frequency (MHz)
	);
	port(
		clk:      in  std_ulogic;
		rst:      in  std_ulogic; -- Active high synchronous reset
		btn:      in  std_ulogic;
		sw:       in  std_ulogic_vector(3 downto 0); -- Slide switches
		data_in:  in  std_ulogic;
		data_drv: out std_ulogic;
		led:      out std_ulogic_vector(3 downto 0); -- LEDs
		stati:out std_logic_vector(4 downto 0)
	);
end entity dht11_sa;

architecture rtl of dht11_sa is

	signal srstn: std_ulogic;
	signal start: std_ulogic;
	signal pe:    std_ulogic;
	signal b:     std_ulogic;
	signal do:    std_ulogic_vector(39 downto 0);
	signal check_parity: std_ulogic;
	signal FSM_stati: std_logic_vector(4 downto 0);

begin
stati <=FSM_stati;
	srstn <= not rst;

	deb: entity work.debouncer(rtl)
	port map(
		clk   => clk,
		srstn => srstn,
		d     => btn,
		q     => open,
		r     => start,
		f     => open,
		a     => open
	);

	u0: entity work.dht11_ctrl(rtl)
	generic map(
		freq => freq
	)
	port map(
		clk      => clk,
		srstn    => srstn,
		start    => start,
		data_in  => data_in,
		data_drv => data_drv,
		pe       => pe,
		b        => b,
		do       => do,
		FSM_stati=>FSM_stati
	);

c_display: entity work.display(rtl)
	generic map( 	N => 4,
			M => 32,
			T => 4)
	port map(
		sw => sw,
		data => do(39 downto 8),
		led => led,
		parity_check => check_parity,
		proto_err => pe,
		busy => b);

c_checksum: entity work.checksum(arc)
  	port map(
	     sresetn => '1',
             data => do,
	     ack => check_parity);

end architecture rtl;

