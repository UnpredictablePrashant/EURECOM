/homes/condemi/Desktop/ds-2017/accumulator/condemi_accumulator.vhd